{# Template for generating RTL pkg addr #}
{# Warn: Keep indentation in phase with module template (cf. addr_snippets) #}
  localparam int {{ofs_name}} = {{ofs_val}};
