{# Template for generating RTL parameter #}          
{# Warn: Keep indentation in phase with module template (cf. param_snippets) #}          
    parameter int {{ default }}
